module cache (
 input [31:0]  address
 ,input read
 ,input write
 ,output [31:0] read_data
 ,output [31:0] write_data 
 
);

 

endmodule
